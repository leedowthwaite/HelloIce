
module Green(input CLK_IN, output GLED5, output RLED1, output RLED2, output RLED3, output RLED4);

	assign GLED5 = 1'b1;

endmodule
